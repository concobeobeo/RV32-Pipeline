module decoder(
	input [31:0] instr,
	output reg stall,
	output reg [1:0] branch_dhazard,
	output reg [1:0] opA,
	output reg [1:0] opB,
	output reg [10:0] data_out);

	// Chu thich:
	// Data_out la ngo ra 11 bits bao gom theo thu tu:
	// {3bit ImmSel, 1bit RegWEn, 4bit ALUSel, 1bit MemRW, 2bit WBSel}
	// Stall tich cuc muc cao
	// opA: 00 rs1, 01 PC, 10 ALU feedback, 11, MEM feedback
	// opB: 00 rs2, 01 Imm, 10 ALU feedback, 11, MEM feedback
	
	reg [4:0] last_rd = 5'bxxxxx;	//buffer cho 2 lenh gan nhat, phuc vu data hazard detect
	reg [4:0] penul_rd = 5'bxxxxx; 	// last of last

	// Define control words 
	// R type instructions
	parameter ADD 	= 9'b000001100;
	parameter SUB 	= 9'b100001100;
	parameter SLL 	= 9'b000101100;
	parameter SLT 	= 9'b001001100;
	parameter SLTU 	= 9'b001101100;
	parameter XOR 	= 9'b010001100;
	parameter SRL 	= 9'b010101100;
	parameter SRA	= 9'b110101100;
	parameter OR 	= 9'b011001100;
	parameter AND	= 9'b011101100;
	// I type instructions
	parameter ADDI 	= 9'b?00000100;
	parameter SLTI 	= 9'b?01000100;
	parameter SLTIU	= 9'b?01100100;
	parameter XORI 	= 9'b?10000100;
	parameter ORI 	= 9'b?11000100;
	parameter ANDI	= 9'b?11100100;
	parameter SLLI 	= 9'b000100100;
	parameter SRLI 	= 9'b010100100;
	parameter SRAI 	= 9'b110100100;
	parameter LW 	= 9'b?01000000;
	// S type instructions
	parameter SW	= 9'b?01001000;
	// B type instructions
	parameter BEQ 	= 9'b?00011000;
	parameter BNE 	= 9'b?00111000;
	parameter BLT 	= 9'b?10011000;
	parameter BLTU	= 9'b?10111000;
	// J type instructions
	parameter JAL  	= 9'b????11011;
	parameter JALR 	= 9'b????11001;
	// U type instructions 
	parameter LUI  	= 9'b????01101;
	parameter AUIPC	= 9'b????00101;


	// 9 bits control.

	wire [10:0] control_word;
	assign control_word = {instr[30], instr[14:12], instr[6:2]};
	always @*
	begin
		casez ({instr[30], instr[14:12], instr[6:2]})
		// R
		ADD: 	data_out = 11'bxxx10000001;
		SUB:	data_out = 11'bxxx10001001;
		SLL:	data_out = 11'bxxx10010001;
		SLT:	data_out = 11'bxxx10011001;
		SLTU:	data_out = 11'bxxx10100001;
		XOR:	data_out = 11'bxxx10101001;
		SRL:	data_out = 11'bxxx10110001;
		SRA:	data_out = 11'bxxx10111001;
		OR: 	data_out = 11'bxxx11000001;
		AND:	data_out = 11'bxxx11001001;
		// 
		ADDI:	data_out = 11'b00010000001;
		SLTI:	data_out = 11'b00010011001;
		SLTIU:	data_out = 11'b00010100001;
		XORI: 	data_out = 11'b00010101001;
		ORI: 	data_out = 11'b00011000001;
		ANDI:	data_out = 11'b00011001001;
		SLLI: 	data_out = 11'b00010010001;
		SRLI: 	data_out = 11'b00010110001;
		SRAI: 	data_out = 11'b00010111001;
		LW:	
			data_out = 11'b00010000000;
		// S
		SW:	data_out = 11'b001000001xx;
		//
		BNE, BEQ, BLT, BLTU: 	
			data_out = 11'b010000000xx;
		// J
		JAL:	data_out = 11'b10010000010;
		JALR:	data_out = 11'b00010000010;
		// 
		LUI:	data_out = 11'b01111011001;
		AUIPC:	data_out = 11'b01110000001; 
		default:data_out = 11'bxxxxxxxxxxx;
		endcase

		// Co rs1, rs2
		// Nhom lenh Branch
		if (instr[6:2] == 5'b11000)
		begin
			// Neu rs1 = rd lenh ke truoc thi opA l� feedback tu tang MEM
			if (instr[19:15]/*rs1*/ == last_rd)
			begin 
				branch_dhazard = 1;
			end
			else if (instr[24:20]/*rs2*/ == last_rd) 
			begin
				branch_dhazard = 2;
			end
			// Neu rs1 hoac rs2 = rd lenh truoc 1 thi opA l� feedback tu tang WB
			/*else if (instr[19:15] == penul_rd)
			begin 
				opA = 2'b11;
				opB = 2'b01;
			end
			else if (instr[24:20] == penul_rd) 
			begin
				opA = 2'b01;
				opB = 2'b11;
			end */ //Do BRANCH O TANG EX NEN KHONG THE BI HAZARD VOI LENH CACH NO 1 LENH
			else 
			begin
				branch_dhazard = 0;
			end
			// cap nhat buffer
			last_rd = 5'bxxxxx;
			penul_rd = 5'bxxxxx;
			stall = 0;
		end
		// Lenh SW
		if (instr[6:2] == 5'b01000)
		begin
			// Neu rs1 = rd lenh ke truoc thi opA l� feedback tu tang MEM
			if (instr[19:15]/*rs1*/ == last_rd)
			begin 
				opA = 2'b10;
				opB = 2'b01;
			end
			else if (instr[24:20]/*rs2*/ == last_rd) 
			begin
				opA = 2'b00;
				opB = 2'b10;
			end
			// Neu rs1 hoac rs2 = rd lenh truoc 1 thi opA l� feedback tu tang WB
			else if (instr[19:15]/*rs1*/ == penul_rd)
			begin 
				opA = 2'b11;
				opB = 2'b01;
			end
			else if (instr[24:20]/*rs2*/ == penul_rd) 
			begin
				opA = 2'b00;
				opB = 2'b11;
			end
			else if (instr[19:15]/*rs1*/ == last_rd && instr[24:20]/*rs2*/ == penul_rd)
			begin
				opA = 2'b10;
				opB = 2'b11;
			end
			else if (instr[19:15]/*rs1*/ == penul_rd && instr[24:20]/*rs2*/ == last_rd)
			begin
				opA = 2'b11;
				opB = 2'b10;
			end
			else 
			begin
				opA = 2'b00;
				opB = 2'b01;
			end
			// cap nhat buffer
			last_rd = 5'bxxxxx;
			penul_rd = 5'bxxxxx;
			stall = 0;
		end
		//-----------------
		// Co rs1, rs2, rd . Nhom lenh R v� 
		else if (instr[6:2] == 5'b01100)
		begin 
			// Neu rs1 hoac rs2 = rd lenh ke truoc thi opA l� feedback tu tang MEM
			if (instr[19:15]/*rs1*/ == last_rd)
			begin 
				opA = 2'b10;
				opB = 2'b00;
			end
			else if (instr[24:20]/*rs2*/ == last_rd)
			begin
				opA = 2'b00;
				opB = 2'b10;
			end
			// Neu rs1 hoac rs2 = rd lenh truoc 1 thi opA l� feedback tu tang WB
			else if (instr[19:15]/*rs1*/ == penul_rd)
			begin 
				opA = 2'b11;
				opB = 2'b00;
			end
			else if (instr[24:20]/*rs2*/ == penul_rd)
			begin
				opA = 2'b00;
				opB = 2'b11;
			end
			else if (instr[19:15]/*rs1*/ == last_rd && instr[24:20]/*rs2*/ == penul_rd)
			begin
				opA = 2'b10;
				opB = 2'b11;
			end
			else if (instr[19:15]/*rs1*/ == penul_rd && instr[24:20]/*rs2*/ == last_rd)
			begin
				opA = 2'b11;
				opB = 2'b10;
			end
			else 
			begin
				opA = 2'b00;
				opB = 2'b00;
			end
			// cap nhat buffer
			penul_rd = last_rd;
			last_rd = instr[11:7];
			stall = 0;
		end 
		// co rs1, rd 
		else if (instr[6:2] == 5'b00000 /*LW*/ || instr[6:2] == 5'b00100 /*IMM*/|| instr[6:2] ==5'b11001 /*JALR*/)
		begin
			// Neu rs1 hoac rs1 = rd lenh ke truoc thi opA l� feedback tu tang MEM
			if (instr[19:15]/*rs1*/ == last_rd)
			begin 
				opA = 2'b10;
				opB = 2'b01;
				if (instr[6:2] == 5'b00000) stall = 1;
			end
			// Neu rs1 hoac rs1 = rd lenh truoc 1 thi opA l� feedback tu tang WB
			else if (instr[19:15]/*rs1*/ == penul_rd)
			begin
				opA = 2'b11;
				opB = 2'b01;
				stall = 0;
			end
			else 
			begin
				opA = 2'b00;
				opB = 2'b01;
				stall = 0;
			end
			// cap nhat buffer
			penul_rd = last_rd;
			last_rd = instr[11:7];
		end
		else begin
			opA = 2'b01;
			opB = 2'b01;
			// cap nhat buffer
			penul_rd = last_rd;
			last_rd = instr[11:7];
			stall = 0;
		end
	end
endmodule 
